library verilog;
use verilog.vl_types.all;
entity tb_change_mode is
end tb_change_mode;
